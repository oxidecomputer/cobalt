// Copyright 2022 Oxide Computer Company
//
// This Source Code Form is subject to the terms of the Mozilla Public
// License, v. 2.0. If a copy of the MPL was not distributed with this
// file, You can obtain one at https://mozilla.org/MPL/2.0/.

package I2C_test;

import I2C::*;

module mkI2cWriteTest (I2cCore);
endmodule: mkI2cWriteTest

endpackage: I2C_test