// This Source Code Form is subject to the terms of the Mozilla Public
// License, v. 2.0. If a copy of the MPL was not distributed with this
// file, You can obtain one at https://mozilla.org/MPL/2.0/.

package LogicSampler;

//
// The LogicSampler package contains primitives to construct a logic sampling
// memory and protocol interface. These primitives allow for the recording of
// typed samples generated by a design (or device I/O pins) and streaming those
// samples somewhere for further analysis.
//

export Offset(..);
export Count(..);
export RecordingHeader(..);
export CommandRequest(..);
export CommandResponse(..);
export Notification(..);
export ControlResponse(..);
export DataResponse(..);

export ControlClient(..);
export ControlServer(..);
export MemoryAddress(..);
export MemoryRequest(..);
export MemoryClient(..);
export MemoryServer(..);

export TriggerFn(..);

export LogicSampler(..);
export LogicSamplingMemory(..);
export ProtocolFrontend(..);

export RequestByte(..);
export ResponseByte(..);
export NotificationByte(..);

export mkLogicSampler;
export mkLogicSamplingBRAM;
export mkByteProtocolFrontend;

import Assert::*;
import BRAM::*;
import ClientServer::*;
import Connectable::*;
import FIFO::*;
import FIFOF::*;
import NumberTypes::*;
import Vector::*;
import StmtFSM::*;


// `Offset` and `Count` types, sized to match a given sample memory depth.
typedef UInt#(TLog#(memory_depth)) Offset#(numeric type memory_depth);
typedef UInt#(TAdd#(TLog#(memory_depth), 1)) Count#(numeric type memory_depth);

//
// Upon playback of a recorded set of samples the sampler provides a header
// indicating the number of samples that where recorded and at what offset in
// the sample stream either the trigger function was matched or the recording
// interrupted.
//
typedef struct {
    Count#(memory_depth) sample_count;
    Offset#(memory_depth) trigger_point_offset;
} RecordingHeader#(numeric type memory_depth) deriving (Bits, Eq, FShow);

//
// `CommandRequest` and `CommandResponse` enums are primitives used in a simple
// control protocol between a protocol frontend and the sampler. There are no
// assumptions made about the latency between a request and response as this is
// implementation dependent.
//
typedef enum {
    Clear,      // Clear the recoding (if any).
    Record,     // Start recording samples.
    Playback,   // Play back recorded samples.
    Stop        // Stop recording or play back of samples.
} CommandRequest deriving (Bits, Eq, FShow);

typedef enum {
    Invalid,    // The command was invalid given the current memory state.
    Ok          // The command was accepted, in progress or completed.
} CommandResponse deriving (Bits, Eq, FShow);

typedef enum {
    TriggerMatch,       // The trigger function was matched.
    RecordingComplete,  // The recording is complete and ready for play back.
    PlaybackComplete    // Play back of the recording has completed.
} Notification deriving (Bits, Eq, FShow);

//
// The `LogicSampler` provides either a `CommandResponse` or `Notification` on a
// given cycle.
//
typedef union tagged {
    CommandResponse Command;
    Notification Notification;
} ControlResponse deriving (Bits, Eq, FShow);

//
// The `LogicSampler` emits either a `RecordingHeader` (at the beginning of play
// back) or a `sample`.
//
typedef union tagged {
    RecordingHeader#(memory_depth) Header;
    sample Sample;
} DataResponse#(numeric type memory_depth, type sample) deriving (Bits, Eq, FShow);

//
// `LogicSampler` control and data Client/Server interfaces.
//
typedef Client#(CommandRequest, ControlResponse) ControlClient;
typedef Server#(CommandRequest, ControlResponse) ControlServer;

//
// Type aliases for the `MemoryClient`/`MemoryServer`, used by the
// `LogicSampler` to store the samples.
//
// Note this should be refactored/made more generic other other types of memory
// are to be supported.
//
typedef BuffIndex#(SizeOf#(Offset#(memory_depth)), memory_depth)
    MemoryAddress#(numeric type memory_depth);

typedef BRAMRequest#(MemoryAddress#(memory_depth), sample)
    MemoryRequest#(numeric type memory_depth, type sample);

typedef BRAMClient#(MemoryAddress#(memory_depth), sample)
    MemoryClient#(numeric type memory_depth, type sample);

typedef BRAM1Port#(MemoryAddress#(memory_depth), sample)
    MemoryServer#(numeric type memory_depth, type sample);

//
// `LogicSampler(..)` implements the sampling and sequencing logic to record and
// play back samples of logic signals. These signals can be either from external
// pins or internal logic.
//
// The `ControlServer` interface is used to issue commands and monitor the state
// of the sampler by listening for notifications. See `mkLogicSampler` for an
// explanation of the control protocol.
//
// The `data` interface is used to stream recorded data from the sampler to a
// client/protocol frontend for processing. This interface is separate from the
// control interface because samples may consists of many bits while control
// primitives are small. This hopefully allows for both paths to only occupy as
// much logic as strictly needed.
//
interface LogicSampler#(numeric type memory_depth, type sample);
    // Sample writer, used to submit samples. Note that this interface is marked
    // always ready since outside logic should under no circumstance be blocked
    // by the sampler nor should it be concerned with whether or not the sampler
    // is ready to receive samples. In case the sampler is unable to record
    // samples they should simply be dropped.
    (* always_ready *) interface Put#(sample) sample;

    // Sampler control and data servers.
    interface ControlServer control;
    interface GetS#(DataResponse#(memory_depth, sample)) data;

    // Sample memory client.
    interface MemoryClient#(memory_depth, sample) memory;
endinterface

// `LogicSamplingMemory` is a trimmed down `LogicSampler` interface which can be
// used when the `LogicSampler` and a memory are instantiated as a single unit.
// See `mkSamplingBRAM` below.
interface LogicSamplingMemory#(numeric type memory_depth, type sample);
    (* always_ready *) interface Put#(sample) sample;
    interface ControlServer control;
    interface GetS#(DataResponse#(memory_depth, sample)) data;
endinterface

//
// Generic protocol frontend interface, which can be connected to some kind of
// bus or protocol interface on one side and a logic sampler on the other.
//
interface ProtocolFrontend#(
        numeric type memory_depth,
        type sample,
        type protocol_request,
        type protocol_response);
    // Protocol frontend.
    interface Server#(protocol_request, protocol_response) protocol;

    // Sample  control/data clients.
    interface ControlClient control;
    interface PutS#(DataResponse#(memory_depth, sample)) data;
endinterface

// Make `ProtocolFrontend` connectable to `LogicSampler`/`LogicSamplingMemory`.
instance Connectable#(
        ProtocolFrontend#(memory_depth, sample, protocol_request, protocol_response),
        LogicSampler#(memory_depth, sample));
    module mkConnection#(
            ProtocolFrontend#(
                memory_depth,
                sample,
                protocol_request,
                protocol_response) frontend,
            LogicSampler#(memory_depth, sample) sampler) (Empty);
        mkConnection(frontend.control, sampler.control);
        mkConnection(frontend.data, sampler.data);
    endmodule
endinstance

instance Connectable#(
        ProtocolFrontend#(memory_depth, sample, protocol_request, protocol_response),
        LogicSamplingMemory#(memory_depth, sample));
    module mkConnection#(
            ProtocolFrontend#(
                memory_depth,
                sample,
                protocol_request,
                protocol_response) frontend,
            LogicSamplingMemory#(memory_depth, sample) memory) (Empty);
        mkConnection(frontend.control, memory.control);
        mkConnection(frontend.data, memory.data);
    endmodule
endinstance

// Trigger function typedef.
typedef (function Bool fn(sample s)) TriggerFn#(type sample);

//
// `mkLogicSampler` instantiates a `LogicSampler` which can be connected to a
// memory in order to implement a `LogicSamplingMemory`. The command protocol
// implemented by this sampler is as follows:
//
// Upon reset the sampler is in its default state, waiting for either a `Record`
// or `Clear` command. Issueing a `Clear` command will reset the sampler state,
// clearing (the metatdata of) a previous recording. Issuing a `Record` command
// starts the sampler causing it to stream samples into memory and applying the
// trigger function to each sample looking for a match. The response to both
// commands is `Ok`, other commands will result in `Invalid`.
//
// While recording samples a `Stop` command can be sent to force the trigger to
// fire and the sampler will respond with `Ok`. Any other command will result in
// `Invalid`.
//
// When the recording is stopped because the trigger function is matched by one
// of the samples the sampler will send a `TriggerMatch` notification. If the
// recording is stopped because a `Stop` command was received no such
// notification will be sent. Upon receiving either a `Stop` command or matching
// the trigger function the sampler will start recording any post trigger sample
// (if configured to do so) and sends a `RecordingComplete` notification when it
// has stopped recording.
//
// At this point the sampler is again in an idle state, waiting for either a
// `Play` or `Clear` command. Issueing a `Clear` command will reset the sampler
// state, clearing (the metatdata of) the recording. Issuing a `Play` command
// will start play back of the recorded data. The response to both commands is
// `Ok`, other commands will result in `Invalid`.
//
// When an `Ok` is received in response to a `Play` command the sampler client
// is expected to use the `data` interface to receive the data. The first item
// received through this interface is a `RecordingHeader` indicating the total
// number of recorded samples as well as the offset in the sample stream where
// the trigger function was matched or the sampler commanded to stop recording.
// After receiving the header the client is expected to `get` the indicated
// number of samples from the `data` interface. Upon sending the last sample the
// sampler indicates the end of play back by sending a `PlaybackComplete`
// notification through the control interface.
//
// Upon completing play back of the recording, the sampler is again in the idle
// state, waiting for either a `Play` or `Clear` command. The recording can be
// played back once more by issuing a `Play` command or cleared by issuing a
// `Clear` command. After clearing the recording the sampler is back in its
// default state and another recording can be started. Note that an explicit
// `Clear` command is required when a recording has completed before a new
// recording can be started.
//
// If the client wishes to stop play back of a recording it can issue a `Stop`
// command during the play back. This will end the play back, clear the data
// interface and the sampler respnds with `Ok` and will return to the idle state
// waiting for either a `Play` or `Clear` command.
//
// The sampler can be tailored to a specific implementation by passing in an
// appropriate trigger function and the desired number of pre/post trigger
// number of samples. Depending on when the trigger function matches or a `Stop`
// command is received the sampler may record a total of `n_samples_pre_trigger
// + n_samples_post_trigger` samples. The sample recorded when either the
// trigger function matched or the recording was stopped is the last sample in
// the pre trigger series.
//
module mkLogicSampler#(
        TriggerFn#(sample) trigger_fn,
        Integer n_samples_pre_trigger,
        Integer n_samples_post_trigger) (LogicSampler#(memory_depth, sample))
            provisos (Bits#(sample, sample_sz));
    staticAssert(n_samples_pre_trigger > 0, "n_samples_pre_trigger == 0");
    staticAssert(
        n_samples_pre_trigger + n_samples_post_trigger <= valueof(memory_depth),
        "n_samples_pre_trigger + n_samples_post_trigger > memory_depth");

    Reg#(SamplerState) state <- mkReg(Clearing);
    RWire#(SamplerState) state_next_request <- mkRWire();

    // Internal rules may need to send control notifications when events occur.
    // They can do so by setting this wire, allowing `do_update_state` to queue
    // a control response.
    RWire#(Notification) sampler_event <- mkRWire();

    // Samples may be wide and/or the trigger function may involve significant
    // combinatorial logic. Since the writer is unaffected by latency as
    // incoming samples can be pipelined, the input is explicitly registered to
    // allow for as much timing slack as possible.
    //
    // The incoming sample FIFO has an unguarded `enq` method, automatically
    // overwriting prior samples if the  is not recording. This satisfies
    // the requirement that samples can always be submitted to the ,
    // irrespective of its state.
    FIFOF#(sample) in_sample <- mkGLFIFOF(True, False);

    // Control/Data I/O.
    FIFO#(CommandRequest) control_request <- mkLFIFO();
    FIFO#(ControlResponse) control_response <- mkSizedFIFO(3);
    FIFO#(DataResponse#(memory_depth, sample)) data_response <- mkFIFO();

    // Writer state.
    Reg#(Count#(memory_depth)) n_samples_recorded <- mkRegU();
    Reg#(Count#(memory_depth)) n_pre_trigger_samples_recorded <- mkRegU();
    Reg#(Count#(memory_depth)) n_post_trigger_samples_recorded <- mkRegU();
    Reg#(Bool) trigger_matched <- mkRegU();

    // Reader state.
    Reg#(Count#(memory_depth)) n_samples_played_back <- mkRegU();

    // Memory client state. The request consists of an address found in one of
    // the counters and an optional incoming sample. Both these pieces are
    // already registered, so the request itself is not explicitly registered.
    // Read responses are registered in `data_response` so no additional
    // register is added here. The memory server may also register its output
    // for one or more cycles, but this is of no consequence to this module
    // other than an additional cycle of latency per sample.
    Reg#(MemoryAddress#(memory_depth)) memory_address <- mkRegU();
    Wire#(MemoryRequest#(memory_depth, sample)) memory_request <- mkWire();
    RWire#(sample) memory_response <- mkRWire();

    Reg#(Bool) memory_request_outstanding <- mkRegU();
    PulseWire memory_request_issued <- mkPulseWire();
    PulseWire memory_response_received <- mkPulseWire();

    function Action set_state(SamplerState state_next) =
        action
            $display("S: ", fshow(state_next));
            state <= state_next;
        endaction;

    function Action complete_request(CommandRequest command, CommandResponse response) =
        action
            $display("R: ", fshow(command), "? ", fshow(response));
            control_response.enq(tagged Command response);
        endaction;

    //
    // Update state if a new state is requested either by internal rules or as a
    // result of control request. Internal state changes have preference over
    // control requests, enforced by the guard on the control request Put
    // interface and the order in the if/else block below.
    //
    (* fire_when_enabled *)
    rule do_state_next (state_next_request.wget matches tagged Valid .state_next);
        set_state(state_next);

        if (sampler_event.wget matches tagged Valid .notification) begin
            $display("N: ", fshow(notification));
            control_response.enq(tagged Notification notification);
        end
    endrule

    (* fire_when_enabled *)
    rule do_control_request (!isValid(state_next_request.wget));
        control_request.deq();

        let request = control_request.first;

        case (tuple2(state, request)) matches
            {AwaitingRecordOrClear, Clear}: begin
                complete_request(request, Ok);
                set_state(Clearing);
            end

            {AwaitingRecordOrClear, Record}: begin
                complete_request(request, Ok);
                set_state(WritingPreTriggerSamples);
            end

            {AwaitingPlaybackOrClear, Clear}: begin
                complete_request(request, Ok);
                set_state(Clearing);
            end

            {AwaitingPlaybackOrClear, Playback}: begin
                complete_request(request, Ok);
                set_state(SendingRecordingHeader);
            end

            default: begin
                complete_request(request, Invalid);
            end
        endcase
    endrule

    //
    // Writer states.
    //

    (* fire_when_enabled *)
    rule do_clear (state == Clearing);
        trigger_matched <= False;
        n_samples_recorded <= 0;
        n_pre_trigger_samples_recorded <= 0;
        n_post_trigger_samples_recorded <= 0;

        in_sample.clear();
        data_response.clear();
        state_next_request.wset(AwaitingRecordOrClear);
    endrule

    (* fire_when_enabled *)
    rule do_record_sample (
            state == WritingPreTriggerSamples ||
            state == WritingPostTriggerSamples);
        // Dequeue the incoming sample and request a write to memory.
        let sample = in_sample.first();
        in_sample.deq();

        memory_request <=
            BRAMRequest{
                write: True,
                responseOnWrite: False,
                address: memory_address,
                datain: sample};

        memory_address <= memory_address + 1;

        // Perform bookkeeping and keep track of the number of recorded samples.
        if (state == WritingPreTriggerSamples) begin
            if (trigger_fn(sample)) begin
                trigger_matched <= True;

                if (n_samples_post_trigger == 0) begin
                    state_next_request.wset(Rewinding);
                    sampler_event.wset(RecordingComplete);
                end
                else begin
                    state_next_request.wset(WritingPostTriggerSamples);
                    sampler_event.wset(TriggerMatch);
                end
            end

            // Clamp the sample counters if the number of pre-trigger samples is
            // reached.
            let saturated = n_pre_trigger_samples_recorded == fromInteger(n_samples_pre_trigger);

            n_pre_trigger_samples_recorded <= n_pre_trigger_samples_recorded + (saturated ? 0 : 1);
            n_samples_recorded <= n_samples_recorded + (saturated ? 0 : 1);
        end
        else if (state == WritingPostTriggerSamples) begin
            n_post_trigger_samples_recorded <= n_post_trigger_samples_recorded + 1;
            n_samples_recorded <= n_samples_recorded + 1;

            if (n_post_trigger_samples_recorded == fromInteger(n_samples_post_trigger - 1)) begin
                state_next_request.wset(Rewinding);
                sampler_event.wset(RecordingComplete);
            end
        end
    endrule

    //
    // Reader states.
    //

    (* fire_when_enabled *)
    rule do_rewind (state == Rewinding);
        //
        // Rewind the sample memory.
        //
        // The `MemoryAddress` and `Count` types are N and N + 1 bits
        // respectively. This allows `Count` to span the entire range of values
        // kept in `MemoryAddress`. Implied in the use of these two types in
        // this module is that a value stored in `Count` never exceeds the
        // maximum value of `MemoryAddress` + 1. Because of this it is safe to
        // truncate the msb of `x`, because in the case this bit is set it means
        // the memory is filled entirely with valid samples and `memory_address`
        // does not need to change. The truncate will cause `x` to be zero in
        // this case.
        //
        // TODO (arjen): determine if one or more asserts can be used to "proof"
        // invariant.
        //
        memory_address <= sbtrctBIUInt(memory_address, truncate(n_samples_recorded));

        n_samples_played_back <= 0;
        memory_request_outstanding <= False;

        data_response.clear();
        state_next_request.wset(AwaitingPlaybackOrClear);
    endrule

    (* fire_when_enabled *)
    rule do_send_playback_header (state == SendingRecordingHeader);
        data_response.enq(
            tagged Header RecordingHeader{
                sample_count: n_samples_recorded,
                trigger_point_offset: truncate(n_pre_trigger_samples_recorded - 1)});

        state_next_request.wset(PlayingBackRecording);
    endrule

    (* fire_when_enabled *)
    rule do_read_memory (
            state == PlayingBackRecording &&
            n_samples_played_back < n_samples_recorded);
        if (!memory_request_outstanding) begin
            memory_request <=
                BRAMRequest{
                    write: False,
                    responseOnWrite: False,
                    address: memory_address,
                    datain: ?};

            memory_request_issued.send();
            memory_address <= memory_address + 1;
        end

        // The `data_response` FIFO automatically provides backpressure by
        // blocking on the `enq` method when samples are not collected.
        if (memory_response.wget matches tagged Valid .sample) begin
            data_response.enq(tagged Sample sample);

            memory_response_received.send();
            n_samples_played_back <= n_samples_played_back + 1;
        end
    endrule

    (* fire_when_enabled *)
    rule do_determine_memory_request_outstanding (state == PlayingBackRecording);
        memory_request_outstanding <=
            (memory_request_outstanding || memory_request_issued) &&
            !memory_response_received;
    endrule

    (* fire_when_enabled *)
    rule do_complete_playback (
            state == PlayingBackRecording &&
            n_samples_played_back == n_samples_recorded);
        sampler_event.wset(PlaybackComplete);
        state_next_request.wset(AwaitingPlaybackOrClear);
    endrule

    //
    // Interfaces.
    //

    interface Put sample = toPut(in_sample);
    interface ControlServer control = toGPServer(control_request, control_response);
    interface GetS data = fifoToGetS(data_response);
    interface MemoryClient memory = toGPClient(memory_request, memory_response);
endmodule: mkLogicSampler

typedef enum {
    Clearing = 0,
    AwaitingRecordOrClear,
    WritingPreTriggerSamples,
    WritingPostTriggerSamples,
    Rewinding,
    AwaitingPlaybackOrClear,
    SendingRecordingHeader,
    PlayingBackRecording
} SamplerState deriving (Bits, Eq, FShow);

//
// `mkSamplingBRAM` combines a `LogicSampler` with a generic BRAM server to make
// a no frils BRAM based logic sampling memory. This is intended for relatively
// small logic sampling applications.
//
module mkLogicSamplingBRAM #(
        TriggerFn#(sample) trigger_fn,
        Integer n_samples_pre_trigger,
        Integer n_samples_post_trigger,
        BRAM_Configure memory_config)
            (LogicSamplingMemory#(memory_depth, sample))
                provisos (Bits#(sample, sample_sz));
    MemoryServer#(memory_depth, sample) memory <- mkBRAM1Server(memory_config);
    LogicSampler#(memory_depth, sample) sampler <-
        mkLogicSampler(
            trigger_fn,
            n_samples_pre_trigger,
            n_samples_post_trigger);

    mkConnection(sampler.memory, memory.portA);

    interface Put sample = sampler.sample;
    interface Control control = sampler.control;
    interface Data data = sampler.data;
endmodule

//
// `mkByteProtocolFrontend` implements a minimal byte oriented protocol frontend
// which can be used to control and stream data from a `LogicSampler` over for
// example a UART, I^2C or SPI interface. The emphasis of this module was to
// test the interfaces of both the `LogicSampler` and `ProtocolFrontend`, so it
// may not be as robust as one would like
//

typedef enum {
    Nop = 32,       // Space
    Interrupt = 73, // I
    Clear = 67,     // C
    Record = 82,    // R
    Playback = 80   // P
} RequestByte deriving (Bits, Eq, FShow);

typedef enum {
    Invalid = 78,   // N
    Ok = 89         // Y
} ResponseByte deriving (Bits, Eq, FShow);

typedef enum {
    TriggerMatch = 84,      // T
    RecordingComplete = 85, // U
    PlaybackComplete = 86   // V
} NotificationByte deriving (Bits, Eq, FShow);

module mkByteProtocolFrontend
        (ProtocolFrontend#(memory_depth, sample, Bit#(8), Bit#(8)))
            provisos (
                Bits#(sample, sample_sz),
                // A sample occupies at most n bytes.
                Div#(sample_sz, 8, n_sample_bytes),
                Add#(sample_sz, a__, TMul#(n_sample_bytes, 8)),
                // The number of sample bytes can be represented by a u32.
                Add#(TLog#(n_sample_bytes), b__, 32),
                // The number of samples can be represented by a u32.
                Add#(SizeOf#(Count#(memory_depth)), c__, 32),
                // The trigger point offset can be represented by a u32.
                Add#(SizeOf#(Offset#(memory_depth)), d__, 32),
                // A counter size which can count max(n_sample_bytes, 4).
                Add#(TLog#(TMax#(n_sample_bytes, 4)), 1, i_sz),
                Add#(n_sample_bytes, e__, TExp#(i_sz)),
                Add#(4, f__, TExp#(i_sz)),
                // SMT magic, bsc wants this in order to compile this module.
                Add#(TMul#(n_sample_bytes, 8), g__, TMul#(TDiv#(TMul#(n_sample_bytes, 8), 8), 8)));
    // Byte protocol server.
    FIFO#(Bit#(8)) in_byte <- mkLFIFO();
    FIFO#(Bit#(8)) out_byte <- mkLFIFO();

    // Sampler control client.
    FIFO#(CommandRequest) sampler_request <- mkFIFO();
    FIFOF#(ControlResponse) sampler_response <- mkLFIFOF();

    // Sample data client.
    Wire#(DataResponse#(memory_depth, sample)) data_response <- mkWire();
    PulseWire data_accepted <- mkPulseWire();

    Reg#(Maybe#(CommandRequest)) request_in_progress <- mkReg(tagged Invalid);
    Reg#(Bool) playback_in_progress <- mkReg(False);

    //
    // Recording serializer.
    //

    Reg#(UInt#(i_sz)) i <- mkRegU();
    Reg#(Count#(memory_depth)) j <- mkRegU();

    function Stmt send_u32(UInt#(32) v) = stream_bytes(out_byte.enq, v, asIfc(i));
    function Stmt send_sample(sample s) = stream_bytes(out_byte.enq, s, asIfc(i));

    FSM playback_seq <- mkFSM(seq
        // Send header, starting with the size of `sample` in bytes.
        send_u32(fromInteger(valueOf(n_sample_bytes)));
        send_u32(extend(data_response.Header.sample_count));
        send_u32(extend(data_response.Header.trigger_point_offset));
        action
            j <= data_response.Header.sample_count;
            data_accepted.send();
        endaction

        // Send the samples.
        while (j > 0) seq
            send_sample(data_response.Sample);
            action
                data_accepted.send();
                j <= j - 1;
            endaction
        endseq
    endseq);

    //
    // Interrupt request handler. This rule runs with pretty much the highest
    // priority and immediately interrupts any in progress playback of a
    // recording. The interrupt is forwarded to the sampler as a `Stop`, forcing
    // a stop if the sampler is recording.
    //
    (* fire_when_enabled *)
    rule do_interrupt (
            !isValid(request_in_progress) &&&
            parse_request(in_byte.first) matches tagged Valid Interrupt);
        in_byte.deq();
        playback_seq.abort();
        request_in_progress <= tagged Valid Stop;
    endrule

    rule do_response (sampler_response.notEmpty && playback_seq.done);
        case (sampler_response.first) matches
            tagged Command .response:
                if (request_in_progress matches tagged Valid .request) begin
                    if (request == Playback && response == Ok) begin
                        playback_seq.start();
                    end

                    out_byte.enq(deparse_response(response));
                    request_in_progress <= tagged Invalid;
                end
                // There does not seem to be a request in progress. Drop the
                // stray response.

            tagged Notification .notification:
                out_byte.enq(deparse_notification(notification));
        endcase

        sampler_response.deq();
    endrule

    (* descending_urgency = "do_interrupt, do_response, do_request" *)
    rule do_request (
            !isValid(request_in_progress) &&
            !sampler_response.notEmpty &&
            playback_seq.done);
        function do_request(r) =
            action
                request_in_progress <= tagged Valid r;
                sampler_request.enq(r);
            endaction;

        if (parse_request(in_byte.first) matches tagged Valid .request) begin
            case (request)
                Nop: out_byte.enq(deparse_response(Ok));
                Interrupt: do_request(Stop);
                Clear: do_request(Clear);
                Record: do_request(Record);
                Playback: do_request(Playback);
            endcase
        end
        else begin
            out_byte.enq(deparse_response(Invalid));
        end

        in_byte.deq();
    endrule

    interface Server protocol = toGPServer(in_byte, out_byte);
    interface ControlClient control = toGPClient(sampler_request, sampler_response);

    interface PutS data;
        method offer = data_response._write;
        method accepted = data_accepted;
    endinterface
endmodule: mkByteProtocolFrontend

//
// ByteProtocolFrontend helpers.
//

function Maybe#(RequestByte) parse_request(Bit#(8) b) =
    case (b)
        32: tagged Valid Nop;
        73: tagged Valid Interrupt;
        67: tagged Valid Clear;
        82: tagged Valid Record;
        80: tagged Valid Playback;
        default: tagged Invalid;
    endcase;

function Bit#(8) deparse_response(CommandResponse r) =
    extend(pack(
        case (r)
            Invalid: ResponseByte'(Invalid);
            Ok: ResponseByte'(Ok);
        endcase));

function Bit#(8) deparse_notification(Notification n) =
    extend(pack(
        case (n)
            TriggerMatch: NotificationByte'(TriggerMatch);
            RecordingComplete: NotificationByte'(RecordingComplete);
            PlaybackComplete: NotificationByte'(PlaybackComplete);
        endcase));

function Vector#(n, Bit#(8)) as_bytes(t v)
        provisos (
            Bits#(t, t_sz),
            Mul#(n, 8, v_sz),
            Add#(t_sz, _, v_sz)) =
    unpack(extend(pack(v)));

function Stmt stream_bytes(function Action a(Bit#(8) b), t v, Reg#(UInt#(i_sz)) i)
        provisos (
            Bits#(t, t_sz),
            Div#(t_sz, 8, n),
            Add#(t_sz, a__, TMul#(n, 8)));
    Vector#(n, Bit#(8)) v_bytes = as_bytes(v);
    return (seq
        for (i <= 0; i < fromInteger(valueOf(n)); i <= i + 1)
            a(v_bytes[i]);
    endseq);
endfunction

endpackage: LogicSampler
