// Copyright 2021 Oxide Computer Company
//
// This Source Code Form is subject to the terms of the Mozilla Public
// License, v. 2.0. If a copy of the MPL was not distributed with this
// file, You can obtain one at https://mozilla.org/MPL/2.0/.

package UART;

export Serializer(..), mkSerializer;
export Deserializer(..), mkDeserializer;
export Serial(..);
export SamplingTransceiver(..), mkSamplingTransceiver;

import Assert::*;
import Connectable::*;
import GetPut::*;
import StmtFSM::*;
import Vector::*;

import BitSampling::*;
import Strobe::*;
import TestUtils::*;


interface Deserializer;
    interface Put#(Bit#(1)) in;
    interface Get#(Bit#(8)) out;
    method Bool waiting_for_start();
    method Bool error();
endinterface

interface Serializer;
    interface Put#(Bit#(8)) in;
    interface Get#(Bit#(1)) out;
endinterface

interface Serial;
    (* prefix = "" *)
    method Action rx((* port = "rx" *) Bit#(1) val);
    method Bit#(1) tx;
endinterface

typedef enum {
    Idle = 0,
    Start,
    Bit0,
    Bit1,
    Bit2,
    Bit3,
    Bit4,
    Bit5,
    Bit6,
    Bit7,
    Stop
} State deriving (Bits, Eq, FShow);

// Cycle through the State enum.
function State next_state(State s) = s == Stop ? Idle : unpack(pack(s) + 1);

module mkSerializer (Serializer);
    Reg#(State) state <- mkReg(Idle);

    // The `in_bits` register holds the current (partial) byte to be shifted out. The Invalid
    // variant indicates a new byte can be clocked in, starting an output bit sequence of a start
    // bit, the byte bits and a stop bit. During this sequence this register will contain the Valid
    // variant and the remaining bits to be shifted out. When a stop bit is shifted out this
    // register is either set to the Invalid variant or the next byte can be clocked in through
    // `in_byte_next`, allowing the bit sequence to restart. The `wset(..)` method of `in_byte_next`
    // is guarded by the Valid bit of `in_byte`. See `Put` interface below.
    //
    // Bit Vectors are used so vector operations are available when shifting bits.
    Reg#(Maybe#(Vector#(8, Bit#(1)))) in_bits <- mkReg(tagged Invalid);
    RWire#(Vector#(8, Bit#(1))) in_byte_next <- mkRWire();

    // Output bit. This register should hold a valid bit at all times. If no more Start, Stop or
    // byte bits are available to shift out this register is set to the Idle bit allowing a
    // downstream consumer to (continue) receive idle bits.
    Reg#(Bit#(1)) out_bit <- mkReg(1); // Idle high.

    // Event generated by the Put interface indicating the pipeline should advance.
    PulseWire shift_out_bit <- mkPulseWire();

    (* no_implicit_conditions, fire_when_enabled *)
    rule do_serialize;
        // Select either the remaining `in_bits` or the next byte if `in_byte_next` is valid.
        // `maybe_in_byte` will be either the Invalid variant, in which case the output bit should
        // be set to idle, or Valid containing some number of bits to be shifted out.
        let maybe_in_bits = isValid(in_byte_next.wget()) ? in_byte_next.wget() : in_bits;

        if (shift_out_bit) begin
            // A bit is being shifted out and a new byte may be clocked in. Determine the next
            // possible states.

            // If next state Idle, in_byte should be empty and output an idle bit.
            let idle = tuple3(Idle, tagged Invalid, 1);

            // If the next state is Start, hold the current bits and output a start bit.
            let start = tuple3(Start, maybe_in_bits, 0);

            // If next state Stop, in_byte should be empty and output a stop bit.
            let stop = tuple3(Stop, tagged Invalid, 1);

            // If the current state is Idle or Stop, the next state can be either Start or Idle
            // depending on whether a new byte is clocked in. Test if `maybe_in_bits` is valid to
            // determine which state to transition to.
            let start_or_idle = isValid(maybe_in_bits) ? start : idle;

            // If shifting bits, keep the tail and output the head. Assume maybe_in_bits is Valid
            // otherwise one of the other states will be selected later.
            let remaining_bits = fromMaybe(?, maybe_in_bits);
            let shift_bit =
                tuple3(
                    next_state(state),
                    // Don't care about the value being shifted in.
                    tagged Valid (shiftOutFrom0(?, remaining_bits, 1)),
                    head(remaining_bits));

            // Select and commit next state.
            match {.state_next, .in_bits_next, .out_bit_next} =
                case (state)
                    Idle: start_or_idle;
                    Bit7: stop;
                    Stop: start_or_idle;
                    default: shift_bit;
                endcase;

            state <= state_next;
            in_bits <= in_bits_next;
            out_bit <= out_bit_next;
        end else begin
            // No bit is shifted out but a new byte may be clocked in so just retain whatever is
            // currently in `maybe_in_bits`.
            in_bits <= maybe_in_bits;
        end
    endrule

    interface Get out;
        method ActionValue#(Bit#(1)) get();
            shift_out_bit.send();
            return out_bit;
        endmethod
    endinterface

    interface Put in;
        method Action put(Bit#(8) d) if (!isValid(in_bits));
            in_byte_next.wset(unpack(d));
        endmethod
    endinterface
endmodule: mkSerializer

(* synthesize *)
module mkSerializerTest (Empty);
    Serializer ser <- mkSerializer();

    mkAutoFSM(seq
        assert_get_eq(ser.out, 1, "expected idle bit");
        assert_get_eq(ser.out, 1, "expected idle bit");
        action
            ser.in.put('h7f);
            assert_get_eq(ser.out, 1, "expected idle bit");
        endaction
        assert_get_eq(ser.out, 0, "expected start bit");
        repeat(7) assert_get_eq(ser.out, 1, "expected high bit");
        assert_get_eq(ser.out, 0, "expected low msb");
        assert_get_eq(ser.out, 1, "expected stop bit");
        assert_get_eq(ser.out, 1, "expected idle bit");
    endseq);

    mkTestWatchdog(15);
endmodule

module mkDeserializer (Deserializer);
    Reg#(State) state <- mkReg(Idle);

    // Next bit received from `Put` interface.
    RWire#(Bit#(1)) in_bit_next <- mkRWire();

    // Bits currently accumulated by the deserializer. The Valid variant holds one or more received
    // bits. The contents of this register are returned upstream via the `Get` interface. A Bit
    // Vector is used here so the shiftInAtX functions can be used.
    Reg#(Maybe#(Vector#(8, Bit#(1)))) out_bits <- mkReg(tagged Invalid);

    // Registered error flag if no Stop bit is received.
    Reg#(Bool) no_stop_bit_received <- mkReg(False);

    // Registered event flag, exposed to upstream to determine if the line is idle and used to guard
    // the `Get` output.
    Reg#(Bool) idle_or_stop <- mkReg(False);

    PulseWire byte_dequeued <- mkPulseWire();

    (* no_implicit_conditions, fire_when_enabled *)
    rule do_deserialize;
        let maybe_out_bits = byte_dequeued ? tagged Invalid : out_bits;

        if (in_bit_next.wget() matches tagged Valid .in_bit) begin
            // A bit is submitted to the deserializer, determine the possible next states.

            // If next state Idle, keep the accumulated bits if upstream has not dequeued, otherwise
            // this will be the Invalid variant.
            let idle = tuple2(Idle, maybe_out_bits);

            // If next state Start, clear the currently accomulated bits.
            let start = tuple2(Start, tagged Valid unpack(0));

            // If next state Stop, keep the currently accumulated bits for upstream to dequeue.
            let stop = tuple2(Stop, maybe_out_bits);

            // If no Stop bit received, clear currently accumulated bits.
            let error = tuple2(Idle, tagged Invalid);

            // While receiving bits, shift bit in msb.
            let accumulated_bits = shiftInAtN(fromMaybe(?, maybe_out_bits), in_bit);
            let receive_bit = tuple2(next_state(state), tagged Valid accumulated_bits);

            // Select and commit next state based on incoming bit.
            match {.state_next, .out_bits_next} =
                case (tuple2(state, in_bit)) matches
                    {Idle, 0}: start;
                    {Idle, 1}: idle;
                    {Bit7, 0}: error;
                    {Bit7, 1}: stop;
                    {Stop, 0}: start;
                    {Stop, 1}: idle;
                    default: receive_bit;
                endcase;

            state <= state_next;
            out_bits <= out_bits_next;

            // Register error strobe.
            no_stop_bit_received <= (state == Bit7 && in_bit == 0);

            // Register Idle or Stop event strobe.
            idle_or_stop <= (state_next == Idle || state_next == Stop);
        end else begin
            // An upstream consumer may have dequeued a byte in which case the Invalid variant
            // should be stored.
            out_bits <= maybe_out_bits;

            // Reset the error strobe so this is a pulse for at most one cycle and can be used to
            // increment a counter.
            no_stop_bit_received <= False;
        end
    endrule

    interface Put in = toPut(in_bit_next);

    interface Get out;
        method ActionValue#(Bit#(8)) get() if (isValid(out_bits) && idle_or_stop);
            byte_dequeued.send();
            return pack(fromMaybe(?, out_bits));
        endmethod
    endinterface

    method error = no_stop_bit_received;
    method waiting_for_start = idle_or_stop;
endmodule: mkDeserializer

(* synthesize *)
module mkSerDesTest (Empty);
    // 10 bit cycles + 2 cycles to latch input/ouput bytes + 1 cycle to assert output.
    mkTestWatchdog(10 + 2 + 1);

    Serializer ser <- mkSerializer();
    Deserializer des <- mkDeserializer();

    mkConnection(ser, des);

    mkAutoFSM(seq
        ser.in.put(8'h55);
        assert_get_eq_display(des.out, 8'h55, "expected 'h55");
    endseq);
endmodule

interface SamplingTransceiver #(numeric type bit_period);
    interface Serial serial;
    interface Put#(Bit#(8)) send;
    interface Get#(Bit#(8)) receive;
    method Bool receive_error();
    method Bool tx_strobe();
endinterface

module mkSamplingTransceiver
        #(Strobe#(any_sz) sample_strobe)
        (SamplingTransceiver#(bit_period))
        provisos (
            Add#(__a, 1, bit_period),         // bit_period > 0.
            Log#(bit_period, bit_period_sz)); // Make bit_period a power of two
    staticAssert(
        2 ** valueof(bit_period_sz) == valueof(bit_period),
        "bit_period should be a power of two");
    staticAssert(valueof(bit_period) > 1, "bit_period should be at least two clock cycles");

    Serializer ser <- mkSerializer();
    Strobe#(bit_period_sz) tx_strobe_ <- mkPowerTwoStrobe(1, 0);

    Deserializer des <- mkDeserializer();
    Strobe#(bit_period_sz) rx_strobe <- mkPowerTwoStrobe(1, 0);
    AsyncBitSampler#(bit_period) rx_sampler <- mkAsyncBitSampler(rx_strobe, NegativePolarity);

    mkConnection(rx_sampler, des);

    (* fire_when_enabled *)
    rule do_tick (sample_strobe);
        rx_strobe.send();
        tx_strobe_.send();
    endrule

    (* fire_when_enabled *)
    rule do_get_next_tx_bit (tx_strobe_);
        let b <- ser.out.get();
    endrule

    interface Serial serial;
        method rx = rx_sampler.in.put;
        method tx = peekGet(ser.out);
    endinterface

    interface Put send = ser.in;
    interface Get receive = des.out;

    method receive_error = des.error;
    method tx_strobe = tx_strobe_._read;
endmodule

// Make Serializer/Deserializer connectable, because we can.
instance Connectable#(Serializer, Deserializer);
    module mkConnection#(Serializer ser, Deserializer des) (Empty);
        mkConnection(ser.out, des.in);
    endmodule
endinstance

instance Connectable#(AsyncBitSampler#(bit_period), Deserializer);
    module mkConnection#(AsyncBitSampler#(bit_period) sampler, Deserializer des) (Empty);
        mkConnection(sampler.out, des.in);

        (* no_implicit_conditions, fire_when_enabled *)
        rule do_search_for_start_bit;
            if (des.waiting_for_start()) begin
                sampler.search_for_bit_edge();
            end
        endrule
    endmodule
endinstance

endpackage : UART
